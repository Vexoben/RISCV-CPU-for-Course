`include "define.v"

module Dispatcher(

);



endmodule