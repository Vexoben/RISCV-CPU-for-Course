`include "define.v"

module Predictor (
   input clk,
   input rst,
   input rdy,
   
);
   
endmodule